module and_gate (
    input       a_i,
    input       b_i,
    output wire c_o
);
  and A1 (c_o, a_i, b_i);
endmodule
