module not_gate (
    input       a_i,
    output wire y_o
);
  not N1 (y_o, a_i);
endmodule