// package fa_package;
//     `include "full_adder.v"
//     `include "add_subtract.v"
// endpackage
