// parameters_pkg.sv
package package_param;

   // Định nghĩa các tham số (parameters)
   parameter RTYPE  = 7'b0110011;
   parameter ITYPE  = 7'b0010011;
   parameter IITYPE = 7'b1100111;
   parameter ILTYPE = 7'b0000011;
   parameter IJTYPE = 7'b1101111;
   parameter STYPE  = 7'b0100011;
   parameter BTYPE  = 7'b1100011;
   parameter U1TYPE = 7'b0110111;
   parameter U2TYPE = 7'b0010111;

endpackage
